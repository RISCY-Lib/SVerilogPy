// Test

module test(
  input logic clk,
  input logic rstz,
  output logic sig
);

endmodule